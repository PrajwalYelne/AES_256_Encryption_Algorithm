module InverseShiftRow(sb,sr);

  input [127:0] sb;
  output [127:0] sr;

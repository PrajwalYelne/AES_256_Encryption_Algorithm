module InverseLastRound(clk,rin,keylastin,fout);
  input clk;
  input [127:0]rin;
  input [127:0]keylastin;
  output [127:0]fout;

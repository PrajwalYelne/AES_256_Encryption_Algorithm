module stupiddeciphertest;

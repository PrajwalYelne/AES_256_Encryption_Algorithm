module MixColumnHelper(rc,mcl);
  input [31:0] rc;
  output [31:0] mcl;

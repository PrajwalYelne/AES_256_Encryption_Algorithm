module InverseSubByte(data,sb);

input [127:0] data;
output [127:0] sb;

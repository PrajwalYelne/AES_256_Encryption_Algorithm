module InverseRounds(clk,data,keyin,rndout);
  input clk;
  input [127:0]data;

module InverseLastRound(clk,rin,keylastin,fout);
  input clk;
  input [127:0]rin;
  

module InverseMixColumn(a,mcl);
  input [127:0] a;
  output [127:0] mcl;
